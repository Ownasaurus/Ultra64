module VHI(output Z);

assign Z = 1'b1;

endmodule
