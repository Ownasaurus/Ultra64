module INVERTED(output Z, input A);

not (Z, A);

endmodule

