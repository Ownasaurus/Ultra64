module AND2(output Z, input A, input B);

and (Z, A, B);

endmodule

