module XOR2(output Z, input A, input B);

xor (Z, A, B);

endmodule

