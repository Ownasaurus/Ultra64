module VLO(output Z);

assign Z = 1'b0;

endmodule
